///////////////////////////////////////////////////////////////////////////////////
// Testbench for Component: OneBitAdder
// Package: FIUSCIS-CDA
// Course: CDA3102 (Computer Architecture), Florida International University
// Developer: Trevor Cickovski
// License: MIT, (C) 2020 All Rights Reserved
///////////////////////////////////////////////////////////////////////////////////

module testbench();
`include "../Test/Test.v"
///////////////////////////////////////////////////////////////////////////////////
// Inputs: A (1-bit)
//         B (1-bit)
//         C (1-bit)
reg A;
reg B;
reg C;
///////////////////////////////////////////////////////////////////////////////////

///////////////////////////////////////////////////////////////////////////////////
// Outputs: S (2-bit)
wire[1:0] S;
///////////////////////////////////////////////////////////////////////////////////

OneBitAdder myAdder(C, A, B, S[0], S[1]);

initial begin
////////////////////////////////////////////////////////////////////////////////////////
// Test: 0+0+0=0 (00)
$display("Testing: 0+0+0=0 (00 in binary)");
A=0; B=0; C=0;  #10; 
verifyEqual2(S, A+B+C);
////////////////////////////////////////////////////////////////////////////////////////

////////////////////////////////////////////////////////////////////////////////////////
// Test: 0+0+1=1 (01)
$display("Testing: 0+0+1=1 (01 in binary)");
A=0; B=0; C=1;  #10; 
verifyEqual2(S, A+B+C);
////////////////////////////////////////////////////////////////////////////////////////

////////////////////////////////////////////////////////////////////////////////////////
// Test: 0+1+0=1 (01)
$display("Testing: 0+1+0=1 (01 in binary)");
A=0; B=1; C=0;  #10; 
verifyEqual2(S, A+B+C);
////////////////////////////////////////////////////////////////////////////////////////

////////////////////////////////////////////////////////////////////////////////////////
// Test: 0+1+1=2 (10)
$display("Testing: 0+1+1=2 (10 in binary)");
A=0; B=1; C=1;  #10; 
verifyEqual2(S, A+B+C);
////////////////////////////////////////////////////////////////////////////////////////

////////////////////////////////////////////////////////////////////////////////////////
// Test: 1+0+0=1 (01)
$display("Testing: 1+0+0=1 (01 in binary)");
A=1; B=0; C=0;  #10; 
verifyEqual2(S, A+B+C);
////////////////////////////////////////////////////////////////////////////////////////

////////////////////////////////////////////////////////////////////////////////////////
// Test: 1+0+1=2 (10)
$display("Testing: 1+0+1=2 (10 in binary)");
A=1; B=0; C=1;  #10; 
verifyEqual2(S, A+B+C);
////////////////////////////////////////////////////////////////////////////////////////

////////////////////////////////////////////////////////////////////////////////////////
// Test: 1+1+0=2 (10)
$display("Testing: 1+1+0=2 (10 in binary)");
A=1; B=1; C=0;  #10; 
verifyEqual2(S, A+B+C);
////////////////////////////////////////////////////////////////////////////////////////

////////////////////////////////////////////////////////////////////////////////////////
// Test: 1+1+1=3 (11)
$display("Testing: 1+1+1=3 (11 in binary)");
A=1; B=1; C=1;  #10; 
verifyEqual2(S, A+B+C);
////////////////////////////////////////////////////////////////////////////////////////


$display("All tests passed.");
end

endmodule

